
module core_x (
);

input  clk;
input  rst_n;
input  struct core_x_in_if;
output struct core_x_out_if;

// feature-1 begin
always @(*) begin
	// detail begin
	// detail end
end
// feature-1 end

endmodule
