
module core_x_sub (
);


endmodule
