
module core_x_cluster ();


endmodule
